library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity char_library is
	port (
			i_clk			: in	std_logic;
			i_rst			: in	std_logic;
			
			i_h_lib_sync	: in	std_logic;
			i_v_lib_sync	: in	std_logic;
			i_sel			: in	integer range 0 to 36;

			o_pix			: out	std_logic
		);
end entity char_library;

architecture RTL of char_library is

	type t_char is array(9 downto 0) of std_logic_vector(0 to 7);
	type t_char_array is array(36 downto 0) of t_char;
	
	constant C_LIB : t_char_array := (
		0 => (	--char = '0'
			0 => "00000000",
			1 => "00111000",
			2 => "01001100",
			3 => "01010100",
			4 => "01100100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
										
		1 => (	--char = '1'
			0 => "00000000",
			1 => "00010000",
			2 => "00110000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		2 => (	--char = '2'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "00000100",
			4 => "00001000",
			5 => "00010000",
			6 => "00100000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),
																			
		3 => (	--char = '3'
			0 => "00000000",
			1 => "01111100",
			2 => "00001000",
			3 => "00010000",
			4 => "00001000",
			5 => "00000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		4 => (	--char = '4'
			0 => "00000000",
			1 => "00001000",
			2 => "00011000",
			3 => "00101000",
			4 => "01001000",
			5 => "01111100",
			6 => "00001000",
			7 => "00001000",
			8 => "00000000",
			9 => "00000000"),	
									
		5 => (	--char = '5'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01111000",
			4 => "00000100",
			5 => "00000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
										
		6 => (	--char = '6'
			0 => "00000000",
			1 => "00011000",
			2 => "00100000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),

		7 => (	--char = '7'
			0 => "00000000",
			1 => "01111100",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "00100000",
			7 => "00100000",
			8 => "00000000",
			9 => "00000000"),
									
		8 => (	--char = '8'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "00111000",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
									
		9 => (	--char = '9'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "00111100",
			5 => "00000100",
			6 => "00001000",
			7 => "00110000",
			8 => "00000000",
			9 => "00000000"),
									
		10 => (	--char = 'A'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01111100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),
									
		11 => (	--char = 'C'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000000",
			4 => "01000000",
			5 => "01000000",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
									
		12 => (	--char = 'D'
			0 => "00000000",
			1 => "01110000",
			2 => "01001000",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01001000",
			7 => "01110000",
			8 => "00000000",
			9 => "00000000"),	
									
		13 => (	--char = 'E'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),
								
		14 => (	--char = 'F'
			0 => "00000000",
			1 => "01111100",
			2 => "01000000",
			3 => "01000000",
			4 => "01111000",
			5 => "01000000",
			6 => "01000000",
			7 => "01000000",
			8 => "00000000",
			9 => "00000000"),	
									
		15 => (	--char = 'G'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000000",
			4 => "01011100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111100",
			8 => "00000000",
			9 => "00000000"),
									
		16 => (	--char = 'H'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01111100",
			5 => "01000100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),
									
		17 => (	--char = 'I'
			0 => "00000000",
			1 => "00111000",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
									
		18 => (	--char = 'L'
			0 => "00000000",
			1 => "01000000",
			2 => "01000000",
			3 => "01000000",
			4 => "01000000",
			5 => "01000000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),
									
		19 => (	--char = 'N'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01100100",
			4 => "01010100",
			5 => "01001100",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),
									
		20 => (	--char = 'O'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
									
		21 => (	--char = 'R'
			0 => "00000000",
			1 => "01111100",
			2 => "01000100",
			3 => "01000100",
			4 => "01111000",
			5 => "01010000",
			6 => "01001000",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),
									
		22 => (	--char = 'S'
			0 => "00000000",
			1 => "00111100",
			2 => "01000000",
			3 => "01000000",
			4 => "00111000",
			5 => "00000100",
			6 => "00000100",
			7 => "01111000",
			8 => "00000000",
			9 => "00000000"),
									
		23 => (	--char = 'T'
			0 => "00000000",
			1 => "01111100",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00010000",
			6 => "00010000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),
									
		24 => (	--char = 'U'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01000100",
			5 => "01000100",
			6 => "01000100",
			7 => "00111000",
			8 => "00000000",
			9 => "00000000"),
									
		25 => (	--char = 'W'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "01010100",
			5 => "01010100",
			6 => "01010100",
			7 => "00101000",
			8 => "00000000",
			9 => "00000000"),
									
		26 => (	--char = 'X'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "00101000",
			4 => "00010000",
			5 => "00101000",
			6 => "01000100",
			7 => "01000100",
			8 => "00000000",
			9 => "00000000"),
									
		27 => (	--char = 'Y'
			0 => "00000000",
			1 => "01000100",
			2 => "01000100",
			3 => "01000100",
			4 => "00101000",
			5 => "00010000",
			6 => "00010000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),
									
		28 => (	--char = 'Z'
			0 => "00000000",
			1 => "01111100",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "01000000",
			7 => "01111100",
			8 => "00000000",
			9 => "00000000"),
									
		29 => (	--char = '?'
			0 => "00000000",
			1 => "00111000",
			2 => "01000100",
			3 => "00000100",
			4 => "00001000",
			5 => "00010000",
			6 => "00000000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),		

		30 => (	--char = '='
			0 => "00000000",
			1 => "00000000",
			2 => "01111100",
			3 => "00000000",
			4 => "01111100",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),	

		31 => (	--char = '+'
			0 => "00000000",
			1 => "00010000",
			2 => "00010000",
			3 => "01111100",
			4 => "00010000",
			5 => "00010000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),										

		32 => (	--char = '-'
			0 => "00000000",
			1 => "00000000",
			2 => "00000000",
			3 => "01111100",
			4 => "00000000",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),	
									
		33 => (	--char = '*'
			0 => "00000000",
			1 => "00000000",
			2 => "01010100",
			3 => "00111000",
			4 => "01111100",
			5 => "00111000",
			6 => "01010100",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),

		34 => (	--char = '/'
			0 => "00000000",
			1 => "00000000",
			2 => "00000100",
			3 => "00001000",
			4 => "00010000",
			5 => "00100000",
			6 => "01000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000"),	
									
		35 => (	--char = '!'
			0 => "00000000",
			1 => "00010000",
			2 => "00010000",
			3 => "00010000",
			4 => "00010000",
			5 => "00000000",
			6 => "00000000",
			7 => "00010000",
			8 => "00000000",
			9 => "00000000"),
									
		36 => (	--char = ' '
			0 => "00000000",
			1 => "00000000",
			2 => "00000000",
			3 => "00000000",
			4 => "00000000",
			5 => "00000000",
			6 => "00000000",
			7 => "00000000",
			8 => "00000000",
			9 => "00000000")
	);

begin

	OUTPUT : process(i_clk, i_rst)
		variable v_H_Pix : integer := 0;
		variable v_V_PIX : integer := 0;
	begin
		if i_rst = '1' then
			v_H_Pix := 0;
			v_V_PIX := 0;
		elsif rising_edge(i_clk) then
			o_pix <= C_LIB(i_sel)(v_V_PIX / 4)(v_H_Pix / 4);
			if i_v_lib_sync = '1' then
				v_H_Pix := 0;
				v_V_PIX := 0;
			elsif i_h_lib_sync = '1' then
				v_H_Pix := 0;
				if v_V_PIX < 39 then
					v_V_PIX := v_V_PIX + 1;
				else
					v_V_PIX := 0;
				end if;
			elsif v_H_Pix < 31 then
				v_H_Pix := v_H_Pix + 1;
			else
				v_H_Pix := 0;
			end if;
		end if;
	end process;
	
end architecture RTL;