LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY char_library IS
	PORT (
			CLK, RST	:	IN		STD_LOGIC;
			SEL		:	IN		INTEGER RANGE 0 TO 27;
			DATA		:	OUT	STD_LOGIC_VECTOR(0 TO 6)
		);
END char_library;

ARCHITECTURE behaviour OF char_library IS
	TYPE char IS ARRAY(8 DOWNTO 0) OF STD_LOGIC_VECTOR(0 TO 6);
	TYPE char_array IS ARRAY(27 DOWNTO 0) OF char;
	
	CONSTANT lib : char_array :=  (
					       0 =>(0 => "0000000",		--char = '0'
									1 => "0011100",
									2 => "0100110",
									3 => "0101010",
									4 => "0110010",
									5 => "0100010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),
										
					       1 =>(0 => "0000000",		--char = '1'
									1 => "0001000",
									2 => "0011000",
									3 => "0001000",
									4 => "0001000",
									5 => "0001000",
									6 => "0001000",
									7 => "0011100",
									8 => "0000000"),

					       2 =>(0 => "0000000",		--char = '2'
									1 => "0011100",
									2 => "0100010",
									3 => "0000010",
									4 => "0000100",
									5 => "0001000",
									6 => "0010000",
									7 => "0111110",
									8 => "0000000"),
																			
					       3 =>(0 => "0000000",		--char = '3'
									1 => "0111110",
									2 => "0000100",
									3 => "0001000",
									4 => "0000100",
									5 => "0000010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),

					       4 =>(0 => "0000000",		--char = '4'
									1 => "0000100",
									2 => "0001100",
									3 => "0010100",
									4 => "0100100",
									5 => "0111110",
									6 => "0000100",
									7 => "0000100",
									8 => "0000000"),	
									
					       5 =>(0 => "0000000",		--char = '5'
									1 => "0111110",
									2 => "0100000",
									3 => "0111100",
									4 => "0000010",
									5 => "0000010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),
										
					      6 => (0 => "0000000",		--char = '6'
									1 => "0001100",
									2 => "0010000",
									3 => "0100000",
									4 => "0111100",
									5 => "0100010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),

					       7 =>(0 => "0000000",		--char = '7'
									1 => "0111110",
									2 => "0000010",
									3 => "0000100",
									4 => "0001000",
									5 => "0010000",
									6 => "0010000",
									7 => "0010000",
									8 => "0000000"),
									
							 8 =>(0 => "0000000",		--char = '8'
									1 => "0011100",
									2 => "0100010",
									3 => "0100010",
									4 => "0011100",
									5 => "0100010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),
									
							 9 =>(0 => "0000000",		--char = '9'
									1 => "0011100",
									2 => "0100010",
									3 => "0100010",
									4 => "0011110",
									5 => "0000010",
									6 => "0000100",
									7 => "0011000",
									8 => "0000000"),
									
							10 =>(0 => "0000000",		--char = 'D'
									1 => "0111000",
									2 => "0100100",
									3 => "0100010",
									4 => "0100010",
									5 => "0100010",
									6 => "0100100",
									7 => "0111000",
									8 => "0000000"),	
									
							11 =>(0 => "0000000",		--char = 'E'
									1 => "0111110",
									2 => "0100000",
									3 => "0100000",
									4 => "0111100",
									5 => "0100000",
									6 => "0100000",
									7 => "0111110",
									8 => "0000000"),
								
							12 =>(0 => "0000000",		--char = 'F'
									1 => "0111110",
									2 => "0100000",
									3 => "0100000",
									4 => "0111100",
									5 => "0100000",
									6 => "0100000",
									7 => "0100000",
									8 => "0000000"),	
									
							13 =>(0 => "0000000",		--char = 'G'
									1 => "0011100",
									2 => "0100010",
									3 => "0100000",
									4 => "0101110",
									5 => "0100010",
									6 => "0100010",
									7 => "0011110",
									8 => "0000000"),
									
							14 =>(0 => "0000000",		--char = 'H'
									1 => "0100010",
									2 => "0100010",
									3 => "0100010",
									4 => "0111110",
									5 => "0100010",
									6 => "0100010",
									7 => "0100010",
									8 => "0000000"),
									
							15 =>(0 => "0000000",		--char = 'L'
									1 => "0100000",
									2 => "0100000",
									3 => "0100000",
									4 => "0100000",
									5 => "0100000",
									6 => "0100000",
									7 => "0111110",
									8 => "0000000"),
									
							16 =>(0 => "0000000",		--char = 'O'
									1 => "0011100",
									2 => "0100010",
									3 => "0100010",
									4 => "0100010",
									5 => "0100010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),
									
							17 =>(0 => "0000000",		--char = 'R'
									1 => "0111110",
									2 => "0100010",
									3 => "0100010",
									4 => "0111100",
									5 => "0101000",
									6 => "0100100",
									7 => "0100010",
									8 => "0000000"),
									
							18 =>(0 => "0000000",		--char = 'T'
									1 => "0111110",
									2 => "0001000",
									3 => "0001000",
									4 => "0001000",
									5 => "0001000",
									6 => "0001000",
									7 => "0001000",
									8 => "0000000"),
									
							19 =>(0 => "0000000",		--char = 'U'
									1 => "0100010",
									2 => "0100010",
									3 => "0100010",
									4 => "0100010",
									5 => "0100010",
									6 => "0100010",
									7 => "0011100",
									8 => "0000000"),
									
							20 =>(0 => "0000000",		--char = 'W'
									1 => "0100010",
									2 => "0100010",
									3 => "0100010",
									4 => "0101010",
									5 => "0101010",
									6 => "0101010",
									7 => "0010100",
									8 => "0000000"),
									
						   21 =>(0 => "0000000",		--char = '?'
									1 => "0011100",
									2 => "0100010",
									3 => "0000010",
									4 => "0000100",
									5 => "0001000",
									6 => "0000000",
									7 => "0001000",
									8 => "0000000"),		

						   22 =>(0 => "0000000",		--char = '='
									1 => "0000000",
									2 => "0111110",
									3 => "0000000",
									4 => "0111110",
									5 => "0000000",
									6 => "0000000",
									7 => "0000000",
									8 => "0000000"),	

						   23 =>(0 => "0000000",		--char = '+'
									1 => "0001000",
									2 => "0001000",
									3 => "0111110",
									4 => "0001000",
									5 => "0001000",
									6 => "0000000",
									7 => "0000000",
									8 => "0000000"),										

						   24 =>(0 => "0000000",		--char = '-'
									1 => "0000000",
									2 => "0000000",
									3 => "0111110",
									4 => "0000000",
									5 => "0000000",
									6 => "0000000",
									7 => "0000000",
									8 => "0000000"),	

							25 =>(0 => "0000000",		--char = '/'
									1 => "0000000",
									2 => "0000010",
									3 => "0000100",
									4 => "0001000",
									5 => "0010000",
									6 => "0100000",
									7 => "0000000",
									8 => "0000000"),								26 =>(0 => "0000000",		--char = '!'
									1 => "0001000",
									2 => "0001000",
									3 => "0001000",
									4 => "0001000",
									5 => "0000000",
									6 => "0000000",
									7 => "0001000",
									8 => "0000000"),
									
							27 =>(0 => "0000000",		--char = ' '
									1 => "0000000",
									2 => "0000000",
									3 => "0000000",
									4 => "0000000",
									5 => "0000000",
									6 => "0000000",
									7 => "0000000",
									8 => "0000000")
								);
BEGIN
	output:PROCESS(CLK, RST)
		VARIABLE count : INTEGER := 0;
	BEGIN
		IF(RST = '1') THEN
			count := 0;
		ELSIF(rising_edge(CLK)) THEN
			IF(count < 9) THEN
				DATA <= lib(SEL)(count);
				count := count + 1;
			ELSE
				DATA <= (OTHERS => '0');
				count := 0;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;