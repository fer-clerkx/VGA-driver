LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY char_library IS
	PORT (
			CLK, RST	:	IN		STD_LOGIC;
			SEL		:	IN		INTEGER RANGE 0 TO 36;
			H_LIB_SYNC : IN STD_LOGIC;
			V_LIB_SYNC : IN STD_LOGIC;
			PIX		:	OUT	STD_LOGIC
		);
END char_library;

ARCHITECTURE behaviour OF char_library IS
	TYPE char IS ARRAY(9 DOWNTO 0) OF STD_LOGIC_VECTOR(0 TO 7);
	TYPE char_array IS ARRAY(36 DOWNTO 0) OF char;
	
	CONSTANT lib : char_array :=  (
					       0 =>(0 => "00000000",		--char = '0'
									1 => "00111000",
									2 => "01001100",
									3 => "01010100",
									4 => "01100100",
									5 => "01000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
										
					       1 =>(0 => "00000000",		--char = '1'
									1 => "00010000",
									2 => "00110000",
									3 => "00010000",
									4 => "00010000",
									5 => "00010000",
									6 => "00010000",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),

					       2 =>(0 => "00000000",		--char = '2'
									1 => "00111000",
									2 => "01000100",
									3 => "00000100",
									4 => "00001000",
									5 => "00010000",
									6 => "00100000",
									7 => "01111100",
									8 => "00000000",
									9 => "00000000"),
																			
					       3 =>(0 => "00000000",		--char = '3'
									1 => "01111100",
									2 => "00001000",
									3 => "00010000",
									4 => "00001000",
									5 => "00000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),

					       4 =>(0 => "00000000",		--char = '4'
									1 => "00001000",
									2 => "00011000",
									3 => "00101000",
									4 => "01001000",
									5 => "01111100",
									6 => "00001000",
									7 => "00001000",
									8 => "00000000",
									9 => "00000000"),	
									
					       5 =>(0 => "00000000",		--char = '5'
									1 => "01111100",
									2 => "01000000",
									3 => "01111000",
									4 => "00000100",
									5 => "00000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
										
					       6 =>(0 => "00000000",		--char = '6'
									1 => "00011000",
									2 => "00100000",
									3 => "01000000",
									4 => "01111000",
									5 => "01000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),

					       7 =>(0 => "00000000",		--char = '7'
									1 => "01111100",
									2 => "00000100",
									3 => "00001000",
									4 => "00010000",
									5 => "00100000",
									6 => "00100000",
									7 => "00100000",
									8 => "00000000",
									9 => "00000000"),
									
							 8 =>(0 => "00000000",		--char = '8'
									1 => "00111000",
									2 => "01000100",
									3 => "01000100",
									4 => "00111000",
									5 => "01000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
									
							 9 =>(0 => "00000000",		--char = '9'
									1 => "00111000",
									2 => "01000100",
									3 => "01000100",
									4 => "00111100",
									5 => "00000100",
									6 => "00001000",
									7 => "00110000",
									8 => "00000000",
									9 => "00000000"),
									
							10 =>(0 => "00000000",		--char = 'A'
									1 => "00111000",
									2 => "01000100",
									3 => "01000100",
									4 => "01000100",
									5 => "01111100",
									6 => "01000100",
									7 => "01000100",
									8 => "00000000",
									9 => "00000000"),
									
							11 =>(0 => "00000000",		--char = 'C'
									1 => "00111000",
									2 => "01000100",
									3 => "01000000",
									4 => "01000000",
									5 => "01000000",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
									
							12 =>(0 => "00000000",		--char = 'D'
									1 => "01110000",
									2 => "01001000",
									3 => "01000100",
									4 => "01000100",
									5 => "01000100",
									6 => "01001000",
									7 => "01110000",
									8 => "00000000",
									9 => "00000000"),	
									
							13 =>(0 => "00000000",		--char = 'E'
									1 => "01111100",
									2 => "01000000",
									3 => "01000000",
									4 => "01111000",
									5 => "01000000",
									6 => "01000000",
									7 => "01111100",
									8 => "00000000",
									9 => "00000000"),
								
							14 =>(0 => "00000000",		--char = 'F'
									1 => "01111100",
									2 => "01000000",
									3 => "01000000",
									4 => "01111000",
									5 => "01000000",
									6 => "01000000",
									7 => "01000000",
									8 => "00000000",
									9 => "00000000"),	
									
							15 =>(0 => "00000000",		--char = 'G'
									1 => "00111000",
									2 => "01000100",
									3 => "01000000",
									4 => "01011100",
									5 => "01000100",
									6 => "01000100",
									7 => "00111100",
									8 => "00000000",
									9 => "00000000"),
									
							16 =>(0 => "00000000",		--char = 'H'
									1 => "01000100",
									2 => "01000100",
									3 => "01000100",
									4 => "01111100",
									5 => "01000100",
									6 => "01000100",
									7 => "01000100",
									8 => "00000000",
									9 => "00000000"),
									
							17 =>(0 => "00000000",		--char = 'I'
									1 => "00111000",
									2 => "00010000",
									3 => "00010000",
									4 => "00010000",
									5 => "00010000",
									6 => "00010000",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
									
							18 =>(0 => "00000000",		--char = 'L'
									1 => "01000000",
									2 => "01000000",
									3 => "01000000",
									4 => "01000000",
									5 => "01000000",
									6 => "01000000",
									7 => "01111100",
									8 => "00000000",
									9 => "00000000"),
									
							19 =>(0 => "00000000",		--char = 'N'
									1 => "01000100",
									2 => "01000100",
									3 => "01100100",
									4 => "01010100",
									5 => "01001100",
									6 => "01000100",
									7 => "01000100",
									8 => "00000000",
									9 => "00000000"),
									
							20 =>(0 => "00000000",		--char = 'O'
									1 => "00111000",
									2 => "01000100",
									3 => "01000100",
									4 => "01000100",
									5 => "01000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
									
							21 =>(0 => "00000000",		--char = 'R'
									1 => "01111100",
									2 => "01000100",
									3 => "01000100",
									4 => "01111000",
									5 => "01010000",
									6 => "01001000",
									7 => "01000100",
									8 => "00000000",
									9 => "00000000"),
									
							22 =>(0 => "00000000",		--char = 'S'
									1 => "00111100",
									2 => "01000000",
									3 => "01000000",
									4 => "00111000",
									5 => "00000100",
									6 => "00000100",
									7 => "01111000",
									8 => "00000000",
									9 => "00000000"),
									
							23 =>(0 => "00000000",		--char = 'T'
									1 => "01111100",
									2 => "00010000",
									3 => "00010000",
									4 => "00010000",
									5 => "00010000",
									6 => "00010000",
									7 => "00010000",
									8 => "00000000",
									9 => "00000000"),
									
							24 =>(0 => "00000000",		--char = 'U'
									1 => "01000100",
									2 => "01000100",
									3 => "01000100",
									4 => "01000100",
									5 => "01000100",
									6 => "01000100",
									7 => "00111000",
									8 => "00000000",
									9 => "00000000"),
									
							25 =>(0 => "00000000",		--char = 'W'
									1 => "01000100",
									2 => "01000100",
									3 => "01000100",
									4 => "01010100",
									5 => "01010100",
									6 => "01010100",
									7 => "00101000",
									8 => "00000000",
									9 => "00000000"),
									
							26 =>(0 => "00000000",		--char = 'X'
									1 => "01000100",
									2 => "01000100",
									3 => "00101000",
									4 => "00010000",
									5 => "00101000",
									6 => "01000100",
									7 => "01000100",
									8 => "00000000",
									9 => "00000000"),
									
							27 =>(0 => "00000000",		--char = 'Y'
									1 => "01000100",
									2 => "01000100",
									3 => "01000100",
									4 => "00101000",
									5 => "00010000",
									6 => "00010000",
									7 => "00010000",
									8 => "00000000",
									9 => "00000000"),
									
							28 =>(0 => "00000000",		--char = 'Z'
									1 => "01111100",
									2 => "00000100",
									3 => "00001000",
									4 => "00010000",
									5 => "00100000",
									6 => "01000000",
									7 => "01111100",
									8 => "00000000",
									9 => "00000000"),
									
						   29 =>(0 => "00000000",		--char = '?'
									1 => "00111000",
									2 => "01000100",
									3 => "00000100",
									4 => "00001000",
									5 => "00010000",
									6 => "00000000",
									7 => "00010000",
									8 => "00000000",
									9 => "00000000"),		

						   30 =>(0 => "00000000",		--char = '='
									1 => "00000000",
									2 => "01111100",
									3 => "00000000",
									4 => "01111100",
									5 => "00000000",
									6 => "00000000",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000"),	

						   31 =>(0 => "00000000",		--char = '+'
									1 => "00010000",
									2 => "00010000",
									3 => "01111100",
									4 => "00010000",
									5 => "00010000",
									6 => "00000000",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000"),										

						   32 =>(0 => "00000000",		--char = '-'
									1 => "00000000",
									2 => "00000000",
									3 => "01111100",
									4 => "00000000",
									5 => "00000000",
									6 => "00000000",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000"),	
									
							33 =>(0 => "00000000",		--char = '*'
									1 => "00000000",
									2 => "01010100",
									3 => "00111000",
									4 => "01111100",
									5 => "00111000",
									6 => "01010100",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000"),

							34 =>(0 => "00000000",		--char = '/'
									1 => "00000000",
									2 => "00000100",
									3 => "00001000",
									4 => "00010000",
									5 => "00100000",
									6 => "01000000",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000"),	
									
							35 =>(0 => "00000000",		--char = '!'
									1 => "00010000",
									2 => "00010000",
									3 => "00010000",
									4 => "00010000",
									5 => "00000000",
									6 => "00000000",
									7 => "00010000",
									8 => "00000000",
									9 => "00000000"),
									
							36 =>(0 => "00000000",		--char = ' '
									1 => "00000000",
									2 => "00000000",
									3 => "00000000",
									4 => "00000000",
									5 => "00000000",
									6 => "00000000",
									7 => "00000000",
									8 => "00000000",
									9 => "00000000")
								);
BEGIN
	output:PROCESS(CLK, RST)
		VARIABLE h_pix : INTEGER := 0;
		VARIABLE v_pix : INTEGER := 0;
	BEGIN
		IF(RST = '1') THEN
			h_pix := 0;
			v_pix := 0;
		ELSIF(rising_edge(CLK)) THEN
			PIX <= lib(SEL)(v_pix / 4)(h_pix / 4);
			IF(V_LIB_SYNC = '1') THEN
				h_pix := 0;
				v_pix := 0;
			ELSIF(H_LIB_SYNC = '1') THEN
				h_pix := 0;
				IF(v_pix < 39) THEN
					v_pix := v_pix + 1;
				ELSE
					v_pix := 0;
				END IF;
			ELSIF(h_pix < 31) THEN
				h_pix := h_pix + 1;
			ELSE
				h_pix := 0;
			END IF;
		END IF;
	END PROCESS;
END ARCHITECTURE;